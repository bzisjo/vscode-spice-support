ADDER - 4 BIT ALL-NAND-GATE BINARY ADDER 
* Example from http://bwrcs.eecs.berkeley.edu/Classes/IcBook/SPICE/Examples/examples.html
*** SUBCIRCUIT DEFINITIONS
.SUBCKT NAND 1 2 3 4 
* NODES: INPUT(2), OUTPUT, VCC 
Q1 9 5 1 QMOD 
D1CLAMP 0 1 DMOD 
Q2 9 5 2 QMOD 
D2CLAMP 0 2 DMOD 
RB 4 5 4K 
R1 4 6 1.6K 
Q3 6 9 8 QMOD 
R2 8 0 1K 
RC 4 7 130 
Q4 7 6 10 QMOD 
DVBEDROP 10 3 DMOD 
Q5 3 8 0 QMOD 
.ENDS NAND

.SUBCKT ONEBIT 1 2 3 4 5 6 
* NODES: INPUT(2), CARRY-IN, OUTPUT, CARRY-OUT, VCC 
X1 1 2 7 6 NAND 
X2 1 7 8 6 NAND 
X3 2 7 9 6 NAND 
X4 8 9 10 6 NAND 
X5 3 10 11 6 NAND 
X6 3 11 12 6 NAND 
X7 10 11 13 6 NAND 
X8 12 13 4 6 NAND 
X9 11 7 5 6 NAND 
.ENDS ONEBIT
.SUBCKT TWOBIT 1 2 3 4 5 6 7 8 9 * NODES: INPUT - BIT0(2) / BIT1(2), OUTPUT - BIT0 / BIT1, * CARRY-IN, CARRY-OUT, VCC 
X1 1 2 7 5 10 9 ONEBIT 
X2 3 4 10 6 8 9 ONEBIT 
.ENDS TWOBIT
.SUBCKT FOURBIT 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 
* NODES: INPUT - BIT0(2) / BIT1(2) / BIT2(2) / BIT3(2), 
* OUTPUT - BIT0 / BIT1 / BIT2 / BIT3, CARRY-IN, 
* CARRY-OUT, VCC 
X1 1 2 3 4 9 10 13 16 15 TWOBIT 
X2 5 6 7 8 11 12 16 14 15 TWOBIT 
.ENDS FOURBIT
*** DEFINE NOMINAL CIRCUIT 
.MODEL DMOD D 
.MODEL QMOD NPN(BF=75 RB=100 CJE=1PF CJC=3PF) 
VCC 99 0 DC 5V 
VIN1A 1 0 PULSE(0 3 0 10NS 10NS 10NS 50NS) 
VIN1B 2 0 PULSE(0 3 0 10NS 10NS 20NS 100NS) 
VIN2A 3 0 PULSE(0 3 0 10NS 10NS 40NS 200NS) 
VIN2B 4 0 PULSE(0 3 0 10NS 10NS 80NS 400NS) 
VIN3A 5 0 PULSE(0 3 0 10NS 10NS 160NS 800NS) 
VIN3B 6 0 PULSE(0 3 0 10NS 10NS 320NS 1600NS) 
VIN4A 7 0 PULSE(0 3 0 10NS 10NS 640NS 3200NS) 
VIN4B 8 0 PULSE(0 3 0 10NS 10NS 1280NS 6400NS) 
X1 1 2 3 4 5 6 7 8 9 10 11 12 0 13 99 FOURBIT RBIT0 9 0 1K 
RBIT1 10 0 1K 
RBIT2 11 0 1K 
RBIT3 12 0 1K 
RCOUT 13 0 1K
*** (FOR THOSE WITH MONEY (AND MEMORY) TO BURN) 
.TRAN 1NS 6400NS 
.END